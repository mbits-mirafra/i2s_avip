`ifndef I2STRANSMITTERSEQUENCEPKG_INCLUDED_
`define I2STRANSMITTERSEQUENCEPKG_INCLUDED_

package I2sTransmitterSequencePkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;
  import I2sTransmitterPkg::*;
  
  `include "I2sTransmitterBaseSeq.sv"

  endpackage : I2sTransmitterSequencePkg
`endif

