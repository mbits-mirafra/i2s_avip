module hvlTop;
 import I2sTestPkg::*;
 import uvm_pkg::*;
 
 initial begin
  run_test("I2sBaseTest");
 end

endmodule : hvlTop

