module hvlTop;
 import I2sTestPkg::*;
 import uvm_pkg::*;
 
 initial begin
  run_test("I2sTest");
 end

endmodule : hvlTop

