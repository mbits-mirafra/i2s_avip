interface I2sInterface;

endinterface
