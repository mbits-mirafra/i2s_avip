`ifndef I2SGLOBALSPKG_INCLUDED_
`define I2SGLOBALSPKG_INCLUDED_

package I2sGlobalsPackage;


typedef enum bit{
    TRUE=1'b1,
    FALSE=1'b0

} hasCoverage_e;


 
endpackage:I2sGlobalsPackage

`endif
