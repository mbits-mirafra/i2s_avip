//--------------------------------------------------------------------------------------------
// HVL_TOP
// It consists of the test_pkg to run the base test
//--------------------------------------------------------------------------------------------
module HvlTop;
 //-------------------------------------------------------
 // Package : Importing Uvm Pakckage and Test Package
 //-------------------------------------------------------
 import I2sTestPkg::*;
 import uvm_pkg::*;
 
 //-------------------------------------------------------
 // run_test for simulation
 //-------------------------------------------------------

 initial begin
  run_test("I2sBaseTest");
 end

endmodule : HvlTop

